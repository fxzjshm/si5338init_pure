import Si5338::*;

module mkTop(Empty);
endmodule
